//New Circuit

module new(N);
output [3:0]N;
assign N = 4'b1010;

endmodule

