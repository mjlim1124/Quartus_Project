module revision(A,B,F);

input A, B;
output F;

//gatelevel(A,B,F);
cassign(A,B,F);
//behav(A,B,F);


endmodule